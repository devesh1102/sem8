// My_Processing_System_tb.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module My_Processing_System_tb (
	);

	wire         my_processing_system_inst_clk_bfm_clk_clk;                       // My_Processing_System_inst_clk_bfm:clk -> [My_Processing_System_inst:clk_clk, My_Processing_System_inst_reset_bfm:clk]
	wire   [3:0] my_processing_system_inst_user_extra_inputs_export;              // My_Processing_System_inst:user_extra_inputs_export -> My_Processing_System_inst_user_extra_inputs_bfm:sig_export
	wire   [3:0] my_processing_system_inst_user_extra_outputs_bfm_conduit_export; // My_Processing_System_inst_user_extra_outputs_bfm:sig_export -> My_Processing_System_inst:user_extra_outputs_export
	wire  [31:0] my_processing_system_inst_user_input_0_export;                   // My_Processing_System_inst:user_input_0_export -> My_Processing_System_inst_user_input_0_bfm:sig_export
	wire  [31:0] my_processing_system_inst_user_input_1_export;                   // My_Processing_System_inst:user_input_1_export -> My_Processing_System_inst_user_input_1_bfm:sig_export
	wire  [31:0] my_processing_system_inst_user_output_bfm_conduit_export;        // My_Processing_System_inst_user_output_bfm:sig_export -> My_Processing_System_inst:user_output_export
	wire         my_processing_system_inst_reset_bfm_reset_reset;                 // My_Processing_System_inst_reset_bfm:reset -> My_Processing_System_inst:reset_reset_n

	My_Processing_System my_processing_system_inst (
		.clk_clk                   (my_processing_system_inst_clk_bfm_clk_clk),                       //                clk.clk
		.reset_reset_n             (my_processing_system_inst_reset_bfm_reset_reset),                 //              reset.reset_n
		.user_extra_inputs_export  (my_processing_system_inst_user_extra_inputs_export),              //  user_extra_inputs.export
		.user_extra_outputs_export (my_processing_system_inst_user_extra_outputs_bfm_conduit_export), // user_extra_outputs.export
		.user_input_0_export       (my_processing_system_inst_user_input_0_export),                   //       user_input_0.export
		.user_input_1_export       (my_processing_system_inst_user_input_1_export),                   //       user_input_1.export
		.user_output_export        (my_processing_system_inst_user_output_bfm_conduit_export)         //        user_output.export
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) my_processing_system_inst_clk_bfm (
		.clk (my_processing_system_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) my_processing_system_inst_reset_bfm (
		.reset (my_processing_system_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (my_processing_system_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_conduit_bfm my_processing_system_inst_user_extra_inputs_bfm (
		.sig_export (my_processing_system_inst_user_extra_inputs_export)  // conduit.export
	);

	altera_conduit_bfm_0002 my_processing_system_inst_user_extra_outputs_bfm (
		.sig_export (my_processing_system_inst_user_extra_outputs_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0003 my_processing_system_inst_user_input_0_bfm (
		.sig_export (my_processing_system_inst_user_input_0_export)  // conduit.export
	);

	altera_conduit_bfm_0003 my_processing_system_inst_user_input_1_bfm (
		.sig_export (my_processing_system_inst_user_input_1_export)  // conduit.export
	);

	altera_conduit_bfm_0004 my_processing_system_inst_user_output_bfm (
		.sig_export (my_processing_system_inst_user_output_bfm_conduit_export)  // conduit.export
	);

endmodule
